---------------------------------------------------------------------------------------------------
-- Author : 
-- Description : 
--   
--   
--   
-- More information (optional) :
--    
--    
---------------------------------------------------------------------------------------------------