package example_package is
 
	constant data_upper_lmt : integer := 15;
	constant data_lower_lmt : integer := 0 ;
 
end package example_package;