library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity generic_reset_bridge_xilinx is
generic (
VENDOR 					: string              := "xilinx"; -- FPGA vendor name, valid values --> "xilinx", "intel", “other”
RESET_ACTIVE_STATUS : std_logic            := '1'; -- '0': active low, '1': active high
SYNCH_FF_NUMBER     : natural range 2 to 5 := 3 -- adjust according to FPGA/SoC family, clock speed and input rate of change
);
port(
	clk 		: in std_logic;
	rst_in 	: in std_logic;
	rst_out	: out std_logic
);
end generic_reset_bridge_xilinx;


architecture behavioral of generic_reset_bridge_xilinx is

signal sync_regs : std_logic_vector(SYNCH_FF_NUMBER -1 downto 0) := (others => (not RESET_ACTIVE_STATUS));
attribute ASYNC_REG : string;
attribute ASYNC_REG of sync_regs : signal is "true";
attribute dont_touch : string;
attribute dont_touch of sync_regs : signal is "true";
attribute iob : string; 
attribute iob of rst_in : port is "true";
begin


	process( clk) begin
		if( rst_in = RESET_ACTIVE_STATUS) then
			sync_regs <= (others => (RESET_ACTIVE_STATUS));
		elsif(rising_Edge(clk)) then
			sync_regs <= sync_regs(SYNCH_FF_NUMBER -2 downto 0) & (not RESET_ACTIVE_STATUS);
		end if;
	end process;
	rst_out <= sync_regs(SYNCH_FF_NUMBER -1 );


end behavioral;