-- to be a self-checking testbench using vhdl report and assert keywords